****************************************
*													*
*			SERIES.CIR							*
*********3 Series X 3 Parallel*************
.include cell_2.lib
.option temp=30
**********First Column************
xcell_01_02 02 01 0201 cell_2 params:area=49  j0=16E-20 j02=1.2E-12
+ jsc=30.5E-3 rs=28e-3 rsh=100000
xcell_02_03 03 02 0302 cell_2 params:area=49  j0=16E-20 j02=1.2E-12
+ jsc=30.5E-3 rs=28e-3 rsh=100000
xcell_03_00 0 03 0003 cell_2 params:area=49  j0=16E-20 j02=1.2E-12
+ jsc=30.5E-3 rs=28e-3 rsh=100000

virrad_01_02  0201  02 dc 900
virrad_02_03  0302  03 dc 900
virrad_03_00  0003  0  dc 900


**********Secondd Column************
xcell_01_12 12 01 1201 cell_2 params:area=49  j0=16E-20 j02=1.2E-12
+ jsc=30.5E-3 rs=28e-3 rsh=100000
xcell_12_13 13 12 1312 cell_2 params:area=49  j0=16E-20 j02=1.2E-12
+ jsc=30.5E-3 rs=28e-3 rsh=100000
xcell_13_00 0  13 0013 cell_2 params:area=49  j0=16E-20 j02=1.2E-12
+ jsc=30.5E-3 rs=28e-3 rsh=100000

virrad_11_12  1201  12 dc 900
virrad_12_13  1312  13 dc 900
virrad_13_00  0013  0  dc 900


**********Third Column**********
xcell_01_22 22 01 2201 cell_2 params:area=49  j0=16E-20 j02=1.2E-12
+ jsc=30.5E-3 rs=28e-3 rsh=100000
xcell_22_23 23 22 2322 cell_2 params:area=49  j0=16E-20 j02=1.2E-12
+ jsc=30.5E-3 rs=28e-3 rsh=100000
xcell_23_00 0  23 0023 cell_2 params:area=49  j0=16E-20 j02=1.2E-12
+ jsc=30.5E-3 rs=28e-3 rsh=100000

virrad_01_22  2201  22 dc 900
virrad_22_23  2322  23 dc 900
virrad_23_00  0023  0 dc 1000



vbias 01 0 dc 0


.plot dc i(vbias)

.dc vbias 0 3.15 0.01
.probe
.end
